//Clock divider 

module clock_div( input wire clk_in, 
						output reg clk_out,
						);
reg counter = 1'b0;
parameter DIVISOR = 						

always @(posedge clk_in)
		begin
		
		end
end module
